`timescale 1ns / 1ps

module glyphs (clk, value, glyph);
	parameter WIDTH = 64;
	parameter ADR_BITS = 6;
	
	input clk;
	input [ADR_BITS-1:0] value;
	output reg [WIDTH-1:0] glyph;
	
	reg [WIDTH-1:0] glyphs [(2**(ADR_BITS+1))-1:0];
	
	initial begin
	
		// To generate other glyphs: http://robojax.com/learn/arduino/8x8LED/
		// NOTE: reverse the order of each row (column: right to left, row: top to bottom)
		glyphs[6'h0] = 64'b0000000000011100001000100010001000100010001000100010001000011100;
		glyphs[6'h1] = 64'b0000000000000100000001000000011000000110000001100000011000000110;
		glyphs[6'h2] = 64'b0000000000001100000100100001000000001000000001000000001000011110;
		glyphs[6'h3] = 64'b0000000000011100001000100010000000011000001000000010001000011100;
		glyphs[6'h4] = 64'b0000000000100010001000100010001000111110001000000010000000100000;
		glyphs[6'h5] = 64'b0000000000111110000000100000001000011110001000000010000000011110;
		glyphs[6'h6] = 64'b0000000000011100000000100000001000011010001001100010001000011100;
		glyphs[6'h7] = 64'b0000000000011110000100000001000000111100000010000000010000000010;
		glyphs[6'h8] = 64'b0000000000011100001000100010001000011100001000100010001000011100;
		glyphs[6'h9] = 64'b0000000000011100001000100010001000111100001000000010001000011100;
		glyphs[6'ha] = 64'b0000000000011000001001000100001001000010011111100100001001000010;
		glyphs[6'hb] = 64'b0000000000011110001000100010001000011110001000100010001000011110;
		glyphs[6'hc] = 64'b0000000000011000001001000000001000000010000000100010010000011000;
		glyphs[6'hd] = 64'b0000000000001110000100100010001000100010001000100001001000001110;
		glyphs[6'he] = 64'b0000000000111110000000100000001000011110000000100000001000111110;
		glyphs[6'hf] = 64'b0000000000111110000000100000001000011110000000100000001000000010;
		glyphs[6'd26] = 64'b0000000000011110001000100010001000011110000000100000001000000000; // P
		glyphs[6'd37] = 64'b0000000000000000000000000100010000101000000100000010100001000100; // x
		glyphs[6'd38] = 64'b0000000000000000000000000000010000000000000001000000000000000000; // :
	
	end
	
	always @(posedge clk)
		glyph <= glyphs[value]; 
	
endmodule

module glyphs2x (clk, value, glyph);
	parameter WIDTH = 4096; // 64x64
	parameter ADR_BITS = 6;
	
	input clk;
	input [ADR_BITS-1:0] value;
	output reg [WIDTH-1:0] glyph;
	
	reg [WIDTH-1:0] glyphs [(2**(ADR_BITS+1))-1:0];
	
	initial begin
		// 0-9
		glyphs[6'h0] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000111111111100001111111110000000000000000000000000000000000000000011111111100000111111111000000000000000000000000000000000000000001111111100000001111111110000000000000000000000000000000000000001111111110000000111111111000000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000011111111100000000111111110000000000000000000000000000000000000001111111110000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111110000000011111111000000000000000000000000000000000000000111111111000000001111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000001111111110000000111111111000000000000000000000000000000000000000011111111000000011111111100000000000000000000000000000000000000001111111110000011111111100000000000000000000000000000000000000000111111111100001111111110000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h1] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111100001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h2] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111110000000011111111110000000000000000000000000000000000000000111100000000000111111111000000000000000000000000000000000000000011000000000000011111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h3] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111100000000011111111110000000000000000000000000000000000000000010000000000000111111111000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000011000000000000001111111110000000000000000000000000000000000000001111100000000001111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h4] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000011111111011111111000000000000000000000000000000000000000000000001111111001111111100000000000000000000000000000000000000000000001111111100111111110000000000000000000000000000000000000000000000111111100011111111000000000000000000000000000000000000000000000111111110001111111100000000000000000000000000000000000000000000111111110000111111110000000000000000000000000000000000000000000011111110000011111111000000000000000000000000000000000000000000011111111000001111111100000000000000000000000000000000000000000011111111000000111111110000000000000000000000000000000000000000001111111000000011111111000000000000000000000000000000000000000001111111100000001111111100000000000000000000000000000000000000000111111100000000111111110000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h5] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111000000000111111111110000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000010000000000000011111111110000000000000000000000000000000000000001111000000000011111111111000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h6] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111110000000011110000000000000000000000000000000000000000011111111110000000000011000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100111111111100000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111110000011111111100000000000000000000000000000000000000011111111110000000111111111000000000000000000000000000000000000001111111111000000011111111100000000000000000000000000000000000000111111111000000000111111110000000000000000000000000000000000000011111111100000000011111111000000000000000000000000000000000000001111111110000000001111111100000000000000000000000000000000000000111111111000000000111111110000000000000000000000000000000000000011111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000001111111110000000111111110000000000000000000000000000000000000000111111111100000111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h7] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h8] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111000001111111110000000000000000000000000000000000000000011111111000000011111111100000000000000000000000000000000000000001111111100000000111111110000000000000000000000000000000000000000111111100000000011111111000000000000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000001111111100000001111111100000000000000000000000000000000000000000111111111000001111111110000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000000111111100000000000000000000000000000000000000011111111000000000011111111000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000001111111111000001111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'h9] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111000001111111110000000000000000000000000000000000000000111111111000000111111111000000000000000000000000000000000000000011111111000000001111111110000000000000000000000000000000000000011111111100000000111111111000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111100000000111111111000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111111000000001111111110000000000000000000000000000000000000001111111110000001111111111000000000000000000000000000000000000000111111111100000111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000111111111110111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000100000000000111111111100000000000000000000000000000000000000000011100000000111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		// A-Z		
		glyphs[6'd10] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000001111111011111111000000000000000000000000000000000000000000000001111111101111111100000000000000000000000000000000000000000000000111111110111111110000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000001111111100111111110000000000000000000000000000000000000000000001111111100011111111000000000000000000000000000000000000000000000111111110001111111100000000000000000000000000000000000000000000011111111000111111111000000000000000000000000000000000000000000011111111100001111111100000000000000000000000000000000000000000001111111100000111111110000000000000000000000000000000000000000000111111110000011111111000000000000000000000000000000000000000000011111111000001111111110000000000000000000000000000000000000000011111111100000111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111110000000000011111111100000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000001111111110000000000001111111100000000000000000000000000000000000111111110000000000000111111111000000000000000000000000000000000111111111000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd11] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111100001111111111111000000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000011111111111110000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111100001111111111111100000000000000000000000000000000000000111111110000000011111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000001111111110000000000000000000000000000000000000111111110000000000111111111000000000000000000000000000000000000011111111000000000011111111100000000000000000000000000000000000001111111100000000001111111110000000000000000000000000000000000000111111110000000000111111111000000000000000000000000000000000000011111111000000000011111111100000000000000000000000000000000000001111111100000000111111111110000000000000000000000000000000000000111111110000111111111111110000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd12] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000011111111111000000011111000000000000000000000000000000000000000001111111111000000000011100000000000000000000000000000000000000000111111111000000000000110000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000001111111110000000000001100000000000000000000000000000000000000000111111111100000000001110000000000000000000000000000000000000000011111111111000000011111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd13] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111100111111111111110000000000000000000000000000000000000000111111110000001111111111100000000000000000000000000000000000000011111111000000011111111110000000000000000000000000000000000000001111111100000000111111111000000000000000000000000000000000000000111111110000000011111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000000111111110000000000000000000000000000000000000011111111000000000011111111000000000000000000000000000000000000001111111100000000001111111100000000000000000000000000000000000000111111110000000000111111110000000000000000000000000000000000000011111111000000000011111111000000000000000000000000000000000000001111111100000000001111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000111111111100000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000000011111111110000000000000000000000000000000000000001111111100000011111111111000000000000000000000000000000000000000111111110011111111111111000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd14] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd15] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd16] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111000000011111000000000000000000000000000000000000000011111111110000000000011100000000000000000000000000000000000000001111111111000000000000110000000000000000000000000000000000000000111111111000000000000001000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000111111111000000111111111111000000000000000000000000000000000000011111111100000011111111111100000000000000000000000000000000000000111111110000001111111111110000000000000000000000000000000000000011111111000000111111111111000000000000000000000000000000000000001111111100000011111111111100000000000000000000000000000000000000111111111000001111111111110000000000000000000000000000000000000011111111100000000001111111000000000000000000000000000000000000001111111110000000000111111100000000000000000000000000000000000000111111111000000000011111110000000000000000000000000000000000000011111111110000000001111111000000000000000000000000000000000000000111111111000000000111111100000000000000000000000000000000000000011111111110000000011111110000000000000000000000000000000000000001111111111000000001111111000000000000000000000000000000000000000011111111111000000111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd17] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000011111111000000000000000000000000000000000000000111111110000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd18] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd19] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011000000000000011111111100000000000000000000000000000000000000001110000000000001111111110000000000000000000000000000000000000000111110000000001111111111000000000000000000000000000000000000000011111100000000111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd20] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000001111111110000000001111111111000000000000000000000000000000000000111111111000000001111111111100000000000000000000000000000000000011111111100000000111111111100000000000000000000000000000000000001111111110000000111111111100000000000000000000000000000000000000111111111000000111111111100000000000000000000000000000000000000011111111100000111111111100000000000000000000000000000000000000001111111110000111111111110000000000000000000000000000000000000000111111111000011111111110000000000000000000000000000000000000000011111111100011111111110000000000000000000000000000000000000000001111111110011111111110000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000011111111101111111111000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111101111111111000000000000000000000000000000000000000000111111111110111111111100000000000000000000000000000000000000000011111111110001111111111000000000000000000000000000000000000000001111111110000111111111100000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000011111111100000111111111100000000000000000000000000000000000000001111111110000001111111111000000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000011111111100000001111111111000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111111000000001111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111111000000000000000000000000000000000000111111111000000000011111111110000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000001111111110000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd21] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd22] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000111111111110000000000000000000000000000000000001111111111000000011111111111000000000000000000000000000000000000111111111100000001111111111100000000000000000000000000000000000011111111111000000111111111110000000000000000000000000000000000001111111111100000111111111111000000000000000000000000000000000000111111111110000011111111111100000000000000000000000000000000000011111111111100001111111111110000000000000000000000000000000000001111111111110001111111111111000000000000000000000000000000000000111111111111000111111111111100000000000000000000000000000000000011111111111100011111111111110000000000000000000000000000000000001111111111111001111111111111000000000000000000000000000000000000111111111111101111111111111100000000000000000000000000000000000011111111111110111111111111110000000000000000000000000000000000001111111111111011111111111111000000000000000000000000000000000000111111101111111111111111111100000000000000000000000000000000000011111110111111111110111111110000000000000000000000000000000000001111111011111111111011111111000000000000000000000000000000000000111111101111111111101111111100000000000000000000000000000000000011111110011111111110111111110000000000000000000000000000000000001111111001111111110011111111000000000000000000000000000000000000111111100111111111001111111100000000000000000000000000000000000011111110011111111100111111110000000000000000000000000000000000001111111000111111110011111111000000000000000000000000000000000000111111100011111110001111111100000000000000000000000000000000000011111110001111111000111111110000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000111111100000000000001111111100000000000000000000000000000000000011111110000000000000111111110000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000111111100000000000001111111100000000000000000000000000000000000011111110000000000000111111110000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000111111100000000000001111111100000000000000000000000000000000000011111110000000000000111111110000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000111111100000000000001111111100000000000000000000000000000000000011111110000000000000111111110000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd23] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111100000000000000000000000000000000000000111111111000000000111111110000000000000000000000000000000000000011111111110000000011111111000000000000000000000000000000000000001111111111000000001111111100000000000000000000000000000000000000111111111100000000111111110000000000000000000000000000000000000011111111111000000011111111000000000000000000000000000000000000001111111111100000001111111100000000000000000000000000000000000000111111111111000000111111110000000000000000000000000000000000000011111111111100000011111111000000000000000000000000000000000000001111111111110000001111111100000000000000000000000000000000000000111111111111100000111111110000000000000000000000000000000000000011111111111110000011111111000000000000000000000000000000000000001111111111111100001111111100000000000000000000000000000000000000111111111111110000111111110000000000000000000000000000000000000011111110111111000011111111000000000000000000000000000000000000001111111011111110001111111100000000000000000000000000000000000000111111101111111000111111110000000000000000000000000000000000000011111110011111100011111111000000000000000000000000000000000000001111111001111111001111111100000000000000000000000000000000000000111111100111111100111111110000000000000000000000000000000000000011111110001111111011111111000000000000000000000000000000000000001111111000111111101111111100000000000000000000000000000000000000111111100001111110111111110000000000000000000000000000000000000011111110000111111111111111000000000000000000000000000000000000001111111000011111111111111100000000000000000000000000000000000000111111100000111111111111110000000000000000000000000000000000000011111110000011111111111111000000000000000000000000000000000000001111111000000111111111111100000000000000000000000000000000000000111111100000011111111111110000000000000000000000000000000000000011111110000001111111111111000000000000000000000000000000000000001111111000000011111111111100000000000000000000000000000000000000111111100000001111111111110000000000000000000000000000000000000011111110000000111111111111000000000000000000000000000000000000001111111000000001111111111100000000000000000000000000000000000000111111100000000111111111110000000000000000000000000000000000000011111110000000001111111111000000000000000000000000000000000000001111111000000000111111111100000000000000000000000000000000000000111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd24] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000111111111100000011111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000011111111110000001111111110000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd25] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000111111110011111111111111100000000000000000000000000000000000000011111111000000011111111110000000000000000000000000000000000000001111111100000000111111111000000000000000000000000000000000000000111111110000000011111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000111111111100000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000000011111111110000000000000000000000000000000000000001111111100111111111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd26] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000111111111100000011111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111110000000011111111100000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000011111111110000001111111110000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd27] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111100011111111111111000000000000000000000000000000000000000111111110000000111111111100000000000000000000000000000000000000011111111000000001111111110000000000000000000000000000000000000001111111100000000111111111000000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111100000000111111111000000000000000000000000000000000000000111111110000000011111111100000000000000000000000000000000000000011111111000000001111111110000000000000000000000000000000000000001111111100000001111111111000000000000000000000000000000000000000111111110001111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000011111111001111111111110000000000000000000000000000000000000000001111111100001111111111000000000000000000000000000000000000000000111111110000011111111110000000000000000000000000000000000000000011111111000000111111111000000000000000000000000000000000000000001111111100000011111111110000000000000000000000000000000000000000111111110000000111111111000000000000000000000000000000000000000011111111000000011111111110000000000000000000000000000000000000001111111100000000111111111000000000000000000000000000000000000000111111110000000011111111110000000000000000000000000000000000000011111111000000000111111111000000000000000000000000000000000000001111111100000000011111111110000000000000000000000000000000000000111111110000000000111111111000000000000000000000000000000000000011111111000000000011111111110000000000000000000000000000000000001111111100000000000111111111000000000000000000000000000000000000111111110000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd28] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111000000001111110000000000000000000000000000000000000000111111111000000000001111000000000000000000000000000000000000000011111111000000000000001100000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000001000000000000000011111111100000000000000000000000000000000000000111000000000000001111111110000000000000000000000000000000000000011111000000000001111111110000000000000000000000000000000000000001111111000000001111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd29] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd30] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000111111111000000001111111110000000000000000000000000000000000000011111111110000001111111111000000000000000000000000000000000000001111111111110011111111111000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd31] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000111111110000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000001111111110000000000011111111100000000000000000000000000000000000011111111000000000001111111110000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000111111110000000001111111110000000000000000000000000000000000000011111111000000000111111110000000000000000000000000000000000000001111111110000000011111111000000000000000000000000000000000000000111111111000000001111111100000000000000000000000000000000000000001111111100000001111111110000000000000000000000000000000000000000111111110000000111111111000000000000000000000000000000000000000011111111000000011111111000000000000000000000000000000000000000001111111110000001111111100000000000000000000000000000000000000000011111111000001111111110000000000000000000000000000000000000000001111111100000111111111000000000000000000000000000000000000000000111111110000011111111000000000000000000000000000000000000000000011111111000001111111100000000000000000000000000000000000000000001111111110000111111110000000000000000000000000000000000000000000011111111000111111111000000000000000000000000000000000000000000001111111100011111111000000000000000000000000000000000000000000000111111110001111111100000000000000000000000000000000000000000000011111111100111111110000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000011111111011111111000000000000000000000000000000000000000000000001111111101111111100000000000000000000000000000000000000000000000111111110111111110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd32] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000001111111100000000000000000000000000000000111111100000000000000000111111110000000000000000000000000000000011111110000000000000000011111111000000000000000000000000000000001111111000000000000000001111111000000000000000000000000000000000111111110000000000000000111111100000000000000000000000000000000011111111000000000000000011111110000000000000000000000000000000001111111100000000000000001111111000000000000000000000000000000000111111110000000000000000111111100000000000000000000000000000000011111111000000000000000011111110000000000000000000000000000000000111111100000000000000011111111000000000000000000000000000000000011111110000111111100001111111100000000000000000000000000000000001111111000011111111000111111110000000000000000000000000000000000111111100011111111100011111110000000000000000000000000000000000011111110001111111110001111111000000000000000000000000000000000001111111100111111111000111111100000000000000000000000000000000000111111110011111111110011111110000000000000000000000000000000000011111111001111111111001111111000000000000000000000000000000000000111111100111111111100111111100000000000000000000000000000000000011111110111111111110011111110000000000000000000000000000000000001111111011111111111001111111000000000000000000000000000000000000111111101111111111110111111100000000000000000000000000000000000011111110111111111111011111100000000000000000000000000000000000001111111011111011111111111110000000000000000000000000000000000000111111111111101111111111111000000000000000000000000000000000000011111111111110111111111111100000000000000000000000000000000000000111111111111001111111111110000000000000000000000000000000000000011111111111100111111111111000000000000000000000000000000000000001111111111100011111111111100000000000000000000000000000000000000111111111110001111111111110000000000000000000000000000000000000011111111111000111111111110000000000000000000000000000000000000001111111111100001111111111000000000000000000000000000000000000000111111111110000111111111100000000000000000000000000000000000000011111111110000011111111110000000000000000000000000000000000000000111111111000001111111111000000000000000000000000000000000000000011111111100000011111111100000000000000000000000000000000000000001111111110000001111111110000000000000000000000000000000000000000111111111000000111111111000000000000000000000000000000000000000011111111000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd33] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000111111111000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000111111111000000000111111111100000000000000000000000000000000000011111111110000000011111111100000000000000000000000000000000000000111111111000000011111111110000000000000000000000000000000000000011111111110000001111111110000000000000000000000000000000000000000111111111000001111111110000000000000000000000000000000000000000001111111110001111111111000000000000000000000000000000000000000000111111111000111111111000000000000000000000000000000000000000000001111111110111111111100000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000001111111111001111111110000000000000000000000000000000000000000000111111111000111111111100000000000000000000000000000000000000000111111111100001111111110000000000000000000000000000000000000000011111111100000111111111100000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000000000011111111110000000111111111100000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000001111111111000000000011111111100000000000000000000000000000000000111111111000000000001111111111000000000000000000000000000000000111111111100000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd34] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000111111111100000000000000000000000000000000111111111100000000000011111111100000000000000000000000000000000001111111110000000000011111111110000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000001111111110000000001111111111000000000000000000000000000000000000111111111100000000111111111000000000000000000000000000000000000001111111110000000111111111100000000000000000000000000000000000000111111111100000011111111100000000000000000000000000000000000000001111111110000011111111110000000000000000000000000000000000000000111111111100001111111110000000000000000000000000000000000000000001111111110001111111111000000000000000000000000000000000000000000111111111100111111111000000000000000000000000000000000000000000001111111110111111111100000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		glyphs[6'd35] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		// x
		glyphs[6'd37] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000011111111111000000000000000000000000000000000000111111111110000001111111111000000000000000000000000000000000000001111111111000001111111111000000000000000000000000000000000000000011111111110000111111111000000000000000000000000000000000000000000111111111000111111111100000000000000000000000000000000000000000011111111110111111111100000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000001111111111001111111110000000000000000000000000000000000000000001111111111000111111111100000000000000000000000000000000000000000111111111100001111111111000000000000000000000000000000000000000111111111100000111111111100000000000000000000000000000000000000111111111100000001111111111000000000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000011111111110000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		// :
		glyphs[6'd38] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		// !
		glyphs[6'd39] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		// shield icon
		glyphs[6'd40] = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	end
	
	always @(posedge clk)
		glyph <= glyphs[value];
		
endmodule
	
